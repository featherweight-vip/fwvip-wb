//----------------------------------------------------------------------
// Created with uvmf_gen version 2023.4
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: This interface performs the fwvip_wb signal monitoring.
//      It is accessed by the uvm fwvip_wb monitor through a virtual
//      interface handle in the fwvip_wb configuration.  It monitors the
//      signals passed in through the port connection named bus of
//      type fwvip_wb_if.
//
//     Input signals from the fwvip_wb_if are assigned to an internal input
//     signal with a _i suffix.  The _i signal should be used for sampling.
//
//     The input signal connections are as follows:
//       bus.signal -> signal_i 
//
//      Interface functions and tasks used by UVM components:
//             monitor(inout TRANS_T txn);
//                   This task receives the transaction, txn, from the
//                   UVM monitor and then populates variables in txn
//                   from values observed on bus activity.  This task
//                   blocks until an operation on the fwvip_wb bus is complete.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
import uvmf_base_pkg_hdl::*;
import fwvip_wb_pkg_hdl::*;
`include "src/fwvip_wb_macros.svh"


interface fwvip_wb_monitor_bfm 
  ( fwvip_wb_if  bus );
  // The pragma below and additional ones in-lined further down are for running this BFM on Veloce
  // pragma attribute fwvip_wb_monitor_bfm partition_interface_xif                                  

`ifndef XRTL
// This code is to aid in debugging parameter mismatches between the BFM and its corresponding agent.
// Enable this debug by setting UVM_VERBOSITY to UVM_DEBUG
// Setting UVM_VERBOSITY to UVM_DEBUG causes all BFM's and all agents to display their parameter settings.
// All of the messages from this feature have a UVM messaging id value of "CFG"
// The transcript or run.log can be parsed to ensure BFM parameter settings match its corresponding agents parameter settings.
import uvm_pkg::*;
`include "uvm_macros.svh"
initial begin : bfm_vs_agent_parameter_debug
  `uvm_info("CFG", 
      $sformatf("The BFM at '%m' has the following parameters: ", ),
      UVM_DEBUG)
end
`endif


  // Structure used to pass transaction data from monitor BFM to monitor class in agent.
`fwvip_wb_MONITOR_STRUCT
  fwvip_wb_monitor_s fwvip_wb_monitor_struct;

  // Structure used to pass configuration data from monitor class to monitor BFM.
 `fwvip_wb_CONFIGURATION_STRUCT
 

  // Config value to determine if this is an initiator or a responder 
  uvmf_initiator_responder_t initiator_responder;
  // Custom configuration variables.  
  // These are set using the configure function which is called during the UVM connect_phase

  tri clock_i;
  tri reset_i;
  tri [31:0] adr_i;
  tri  cyc_i;
  tri  ack_i;
  tri  err_i;
  tri [3:0] sel_i;
  tri  stb_i;
  tri  we_i;
  tri [31:0] dat_w_i;
  tri [31:0] dat_r_i;
  assign clock_i = bus.clock;
  assign reset_i = bus.reset;
  assign adr_i = bus.adr;
  assign cyc_i = bus.cyc;
  assign ack_i = bus.ack;
  assign err_i = bus.err;
  assign sel_i = bus.sel;
  assign stb_i = bus.stb;
  assign we_i = bus.we;
  assign dat_w_i = bus.dat_w;
  assign dat_r_i = bus.dat_r;

  // Proxy handle to UVM monitor
  fwvip_wb_pkg::fwvip_wb_monitor  proxy;
  // pragma tbx oneway proxy.notify_transaction                 

  // pragma uvmf custom interface_item_additional begin
  // pragma uvmf custom interface_item_additional end
  
  //******************************************************************                         
  task wait_for_reset();// pragma tbx xtf  
    @(posedge clock_i) ;                                                                    
    do_wait_for_reset();                                                                   
  endtask                                                                                   

  // ****************************************************************************              
  task do_wait_for_reset(); 
  // pragma uvmf custom reset_condition begin
    wait ( reset_i === 1 ) ;                                                              
    @(posedge clock_i) ;                                                                    
  // pragma uvmf custom reset_condition end                                                                
  endtask    

  //******************************************************************                         
 
  task wait_for_num_clocks(input int unsigned count); // pragma tbx xtf 
    @(posedge clock_i);  
                                                                   
    repeat (count-1) @(posedge clock_i);                                                    
  endtask      

  //******************************************************************                         
  event go;                                                                                 
  function void start_monitoring();// pragma tbx xtf    
    -> go;
  endfunction                                                                               
  
  // ****************************************************************************              
  initial begin                                                                             
    @go;                                                                                   
    forever begin                                                                        
      @(posedge clock_i);  
      do_monitor( fwvip_wb_monitor_struct );
                                                                 
 
      proxy.notify_transaction( fwvip_wb_monitor_struct );
 
    end                                                                                    
  end                                                                                       

  //******************************************************************
  // The configure() function is used to pass agent configuration
  // variables to the monitor BFM.  It is called by the monitor within
  // the agent at the beginning of the simulation.  It may be called 
  // during the simulation if agent configuration variables are updated
  // and the monitor BFM needs to be aware of the new configuration 
  // variables.
  //
    function void configure(fwvip_wb_configuration_s fwvip_wb_configuration_arg); // pragma tbx xtf  
    initiator_responder = fwvip_wb_configuration_arg.initiator_responder;
  // pragma uvmf custom configure begin
  // pragma uvmf custom configure end
  endfunction   


  // ****************************************************************************  
            
  task do_monitor(output fwvip_wb_monitor_s fwvip_wb_monitor_struct);
    //
    // Available struct members:
    //     //    fwvip_wb_monitor_struct.adr
    //     //    fwvip_wb_monitor_struct.dat
    //     //    fwvip_wb_monitor_struct.sel
    //     //    fwvip_wb_monitor_struct.we
    //     //
    // Reference code;
    //    How to wait for signal value
    //      while (control_signal === 1'b1) @(posedge clock_i);
    //    
    //    How to assign a struct member, named xyz, from a signal.   
    //    All available input signals listed.
    //      fwvip_wb_monitor_struct.xyz = adr_i;  //    [31:0] 
    //      fwvip_wb_monitor_struct.xyz = cyc_i;  //     
    //      fwvip_wb_monitor_struct.xyz = ack_i;  //     
    //      fwvip_wb_monitor_struct.xyz = err_i;  //     
    //      fwvip_wb_monitor_struct.xyz = sel_i;  //    [3:0] 
    //      fwvip_wb_monitor_struct.xyz = stb_i;  //     
    //      fwvip_wb_monitor_struct.xyz = we_i;  //     
    //      fwvip_wb_monitor_struct.xyz = dat_w_i;  //    [31:0] 
    //      fwvip_wb_monitor_struct.xyz = dat_r_i;  //    [31:0] 
    // pragma uvmf custom do_monitor begin
    // UVMF_CHANGE_ME : Implement protocol monitoring.  The commented reference code 
    // below are examples of how to capture signal values and assign them to 
    // structure members.  All available input signals are listed.  The 'while' 
    // code example shows how to wait for a synchronous flow control signal.  This
    // task should return when a complete transfer has been observed.  Once this task is
    // exited with captured values, it is then called again to wait for and observe 
    // the next transfer. One clock cycle is consumed between calls to do_monitor.
    while (cyc_i !== 1'b1 || stb_i !== 1'b1 || ack_i !== 1'b1) begin
        @(posedge clock_i);
    end
    fwvip_wb_monitor_struct.adr = adr_i;
    if (we_i) begin
        fwvip_wb_monitor_struct.dat = dat_w_i;
    end else begin
        fwvip_wb_monitor_struct.dat = dat_r_i;
    end
    fwvip_wb_monitor_struct.sel = sel_i;
    fwvip_wb_monitor_struct.we = we_i;

    // pragma uvmf custom do_monitor end
  endtask         
  
 
endinterface

// pragma uvmf custom external begin
// pragma uvmf custom external end

