
`include "uvm_macros.svh"
package fwvip_wb_tests_pkg;
    import uvm_pkg::*;
    import fwvip_wb_env_pkg::*;
    import fwvip_wb_pkg::*;

    `include "fwvip_wb_test_base.svh"
    `include "fwvip_wb_test_init.svh"

endpackage

