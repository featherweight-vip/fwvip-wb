
package fwvip_wb_bfm_pkg;
    parameter int ADDR_WIDTH_MAX = 64;
    parameter int DATA_WIDTH_MAX = 64;

endpackage
